`define CORDIC_NTAB 16
`define M_PI        3.141592653589793
`define K           1.646760258121066
`define CORDIC_1K   32'h000026dd   
`define PI          32'h0000c90f
`define TWO_PI      32'h0001921f 
`define HALF_PI     32'h00006487

`define NEG_PI      32'hffff36f1
`define NEG_TWO_PI  32'hfffe6de1
`define NEG_HALF_PI 32'hffff9b79
`define NEG_CORDIC_1K 32'hffffd923

// integer bits are 31:14