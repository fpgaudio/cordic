module cordic

endmodule