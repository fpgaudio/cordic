`ifndef __GLOBALS__
`define __GLOBALS__

// UVM Globals
localparam P_FIXED_NAME = "../rad.txt";
localparam SIN_OUT_NAME = "../sin_out.txt";
localparam SIN_CMP_NAME = "../sin.txt";
localparam COS_OUT_NAME = "../cos_out.txt";
localparam COS_CMP_NAME = "../cos.txt";


localparam CLOCK_PERIOD = 10;

`endif
 